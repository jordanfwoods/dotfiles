-------------------------------------
-- Originator       : Jordan Woods --
-- Last Modified By : Jordan Woods --
-- Last Modified    : <>/<>/<>     --
-------------------------------------
--
--------------------------------------------------------------------------------
-- <Module Name>.sv = <Basic Description>                                     --
-- This module does the following:                                            --
-- 1) TBD                                                                     --
--                                                                            --
-- Revision History                                                           --
-- <>/<>/<> - JFW - Initial Release                                           --
--------------------------------------------------------------------------------
--
------------------------------------------------------------
-- Copyright 2021, Space Micro, Inc. All rights reserved. --
------------------------------------------------------------
