b_example : block
begin
   q <= d when a = '1' else '0';
end block;
