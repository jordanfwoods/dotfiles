----------------------------------------------
-- Originator       : Jordan Woods          --
-- Last Modified By : $Author::           $ --
-- Last Modified    : $Date::             $ --
-- SVN Revision     : $Rev::              $ --
----------------------------------------------
--
--------------------------------------------------------------------------------
-- <Module Name> = <Basic Description>                                        --
-- This module does the following:                                            --
-- 1) TBD                                                                     --
--                                                                            --
-- Revision History                                                           --
-- <>/<>/<> - JFW - Initial Release                                           --
--------------------------------------------------------------------------------
--
------------------------------------------------------------
-- Copyright 2022, Space Micro, Inc. All rights reserved. --
------------------------------------------------------------
