out1 <= in1 or in2;
out2 <= in1 nor in2;
out3 <= in1 and in2;
out4 <= in1 nand in2;
out5 <= in1 xor in2;
out6 <= in1 xnor in2;
out7 <= not in1;
