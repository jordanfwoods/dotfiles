for ID in range loop
    {sequential statement}
end loop;
