--------------------------------------------------------------------------------
-- REPLACE_BY_PROJECT
--------------------------------------------------------------------------------
--
-- Filename          : REPLACE_BY_FUNCTION.vhd
-- VHDL Entity       : REPLACE_BY_FUNCTION
--      Architecture : rtl/behave
--      Library      : REPLACE_BY_PROJECT
--
-- Created:
--          by - REPLACE_BY_NAME
--          at - REPLACE_BY_DATE_YYYY_MM_DD
--
--------------------------------------------------------------------------------
-- Copyright (c) 2023, ASML
--------------------------------------------------------------------------------
-- Purpose      :
--
--------------------------------------------------------------------------------
-- Comment      :
--
--------------------------------------------------------------------------------
-- Assumptions  :
--
--------------------------------------------------------------------------------
-- Limitations  :
--
--------------------------------------------------------------------------------
-- Known Errors :
--
--------------------------------------------------------------------------------
-- Specification Reference :
--
--------------------------------------------------------------------------------
-- History:
-- Date         Author                  Comment
-- REPLACE_BY_DATE_YYYY_MM_DD   REPLACE_BY_NAME      Initial design
--
--
--------------------------------------------------------------------------------
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity REPLACE_BY_FUNCTION is
end entity REPLACE_BY_FUNCTION;

architecture rtl of REPLACE_BY_FUNCTION is
begin
end architecture rtl;
