//////////////////////////////////////////////
// Originator       : Jordan Woods          //
// Last Modified By : $Author::           $ //
// Last Modified    : $Date::             $ //
// SVN Revision     : $Rev::              $ //
//////////////////////////////////////////////
//
////////////////////////////////////////////////////////////////////////////////
// <Module Name> = <Basic Description>                                        //
// This module does the following:                                            //
// 1) TBD                                                                     //
//                                                                            //
// Manual Revision History                                                    //
// <>/<>/<> - JFW - Initial Release                                           //
////////////////////////////////////////////////////////////////////////////////
//
////////////////////////////////////////////////////////////
// Copyright 2021, Space Micro, Inc. All rights reserved. //
////////////////////////////////////////////////////////////
