----------------------------------------------
-- Originator       : Jordan Woods          --
-- Last Modified By : $Author::           $ --
-- Last Modified    : $Date::             $ --
-- SVN Revision     : $Rev::              $ --
----------------------------------------------
--
--------------------------------------------------------------------------------
-- <Module Name> = <Basic Description>                                        --
-- This module does the following:                                            --
-- 1) TBD                                                                     --
--                                                                            --
-- Revision History                                                           --
-- <>/<>/<> - JFW - Initial Release                                           --
--------------------------------------------------------------------------------
--
------------------------------------------------------------
-- Copyright 2023, Space Micro, Inc. All rights reserved. --
------------------------------------------------------------

  ----------------
  -- Parameters --
  ----------------

  ------------------------
  -- Signal Definitions --
  ------------------------

  -------------
  -- Aliases --
  -------------

  ------------------------------
  -- Component Instantiations --
  ------------------------------

  -------------------------
  -- Combinatorial logic --
  -------------------------

  ----------------------
  -- Sequential logic --
  ----------------------

