function bypass(inp: std_logic) return std_logic is
begin
   return inp;
end bypass;
