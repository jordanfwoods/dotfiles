package example_package is
   procedure print(active: boolean);
   type ABC is (A, B, C);
end example_package;
