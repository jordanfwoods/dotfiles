package body example_package is
   procedure print(active: boolean) is
   begin
      if active then
         -- do something
      end if;
   end print;
end example_package;
