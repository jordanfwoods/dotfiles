procedure bypass2(inp: in std_logic; outp: inout std_logic)is
begin
  outp <= inp;
end bypass2;
