architecture rtl of example_entity is
   -- Put your signal/type declarations here
   signal output : std_logic;
   variable v_cnt : integer;
begin
   -- Put your assignments here
   your_output0 <= your_input0;
   your_output1 <= your_input1;

   -- Put your instantiations here

   -- Put your processes here
end rtl;
