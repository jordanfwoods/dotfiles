if expr1 then
   counter <= 0;
elsif expr2 then
   counter <= 1;
else
   counter <= 2;
endif;
