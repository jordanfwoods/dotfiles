while expr loop
   {sequential statement}
end loop;
