case counter is
   when 0 => {sequential statement}
   when 1 => {sequential statement}
   when others => null;
end case;
